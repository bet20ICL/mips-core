module JR_tb();



endmodule