module ALU();

endmodule