module testbench();

endmodule