module lw_harvard_tb();



endmodule