module instruction_ram (
    input logic clk
);
    
endmodule