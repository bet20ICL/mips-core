module convert_endian(
    input logic[31:0] in;
    output logic[31:0] out;
);

    

endmodule 