module lw_harvard_tb.v();

err

endmodule