module regfile(
    input logic[]
);

endmodule