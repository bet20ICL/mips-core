module alu_control(
    input logic[5:0] alu_opcode,
    input logic[5:0] alu_fcode,
    output logic[2:0] alu_control_out
);

endmodule