module data_ram (
    input logic clk
);
    
endmodule