//Combinatorial read of data, no write

module instruction_ram (
    input logic[31:0]  instr_address,
    output logic[31:0]   instr_readdata
);
    
endmodule